library ieee;
use ieee.std_logic_1164.all;

package utility_pkg is

  type std_logic_vector_array_t is array (natural range <>) of std_logic_vector;
  type std_logic_vector_array_3D_t is array (natural range <>) of std_logic_vector_array_t;

end package utility_pkg;

package body utility_pkg is
end package body utility_pkg;
