library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.gt_pkg.all;
use work.axi_lane_pkg.all;


entity AXI_interface is
    port( 
        eth_gtrefclk_p : in std_logic;
        eth_gtrefclk_n : in std_logic;
        -- Ethernet SFP lane
        txn_eth_sfp : out std_logic;
        txp_eth_sfp : out std_logic;
        rxn_eth_sfp : in  std_logic;
        rxp_eth_sfp : in  std_logic;
        
        -- Ethernet addresses selection (group1 [1, Tx], group2 [2, Rx] or VIO [0])
        eth_addr_sel : in std_logic_vector(1 downto 0);
        
        -- IIC
        sda : inout std_logic;
        scl : inout std_logic;
        
        -- synch and shared data
        clk_sys  : in  std_logic;
        rxusrclk : in  std_logic;
        txusrclk : in  std_logic;
        to_axi   : in  to_axi_t;
        from_axi : out from_axi_t
    );
end AXI_interface;

architecture Behavioral of AXI_interface is

    -- AXI MM Interface
    signal resetn_axi    : std_logic; -- generated by the AXI master signal
    
    signal m_axi_lane_awaddr  : axi_lane_awaddr_t;
    signal m_axi_lane_awvalid : axi_lane_awvalid_t;
    signal m_axi_lane_awready : axi_lane_awready_t := (others => '0');
    signal m_axi_lane_wdata   : axi_lane_wdata_t;
    signal m_axi_lane_wstrb   : axi_lane_wstrb_t;
    signal m_axi_lane_wvalid  : axi_lane_wvalid_t;
    signal m_axi_lane_wready  : axi_lane_wready_t := (others => '0');
    signal m_axi_lane_bresp   : axi_lane_bresp_t := (others => (others => '0'));
    signal m_axi_lane_bvalid  : axi_lane_bvalid_t := (others => '0');
    signal m_axi_lane_bready  : axi_lane_bready_t;
    signal m_axi_lane_araddr  : axi_lane_araddr_t;
    signal m_axi_lane_arvalid : axi_lane_arvalid_t;
    signal m_axi_lane_arready : axi_lane_arready_t := (others => '0');
    signal m_axi_lane_rdata   : axi_lane_rdata_t := (others => (others => '0'));
    signal m_axi_lane_rresp   : axi_lane_rresp_t := (others => (others => '0'));
    signal m_axi_lane_rvalid  : axi_lane_rvalid_t := (others => '0');
    signal m_axi_lane_rready  : axi_lane_rready_t;
    
    signal m_axi_aux_awaddr  : std_logic_vector(31 downto 0);
    signal m_axi_aux_awvalid : std_logic;
    signal m_axi_aux_awready : std_logic;
    signal m_axi_aux_wdata   : std_logic_vector(31 downto 0);
    signal m_axi_aux_wstrb   : std_logic_vector(3 downto 0);
    signal m_axi_aux_wvalid  : std_logic;
    signal m_axi_aux_wready  : std_logic;
    signal m_axi_aux_bresp   : std_logic_vector(1 downto 0);
    signal m_axi_aux_bvalid  : std_logic;
    signal m_axi_aux_bready  : std_logic;
    signal m_axi_aux_araddr  : std_logic_vector(31 downto 0);
    signal m_axi_aux_arvalid : std_logic;
    signal m_axi_aux_arready : std_logic;
    signal m_axi_aux_rdata   : std_logic_vector(31 downto 0);
    signal m_axi_aux_rresp   : std_logic_vector(1 downto 0);
    signal m_axi_aux_rvalid  : std_logic;
    signal m_axi_aux_rready  : std_logic;
    
    signal axi_gpio_state        : std_logic_vector(31 downto 0);
    signal axi_gpio_state_asynch : std_logic_vector(31 downto 0);
    
    signal axi_gpio_ctrl_async   : std_logic_vector(11 downto 0); -- := "00000000 0100"; -- := "10101010 0100";
    signal axi_gpio_ctrl         : std_logic_vector(3 downto 0); -- := "0100";

begin

    axi_gpio_state_asynch <= to_axi.slide_count(6 downto 0) & to_axi.lol_count & to_axi.lol_ovf & to_axi.odds_count(4 downto 0) & to_axi.temp & to_axi.ready; -- 7 + 8 + 1 + 5 + 10 + 1 bits

    bus_synch_rx_to_axi: entity work.bus_synch
      generic map ( NBITS => 32 ) 
      port map (
        clk            => clk_sys,
        clk_start      => rxusrclk,
        data_asynch_in => axi_gpio_state_asynch, 
        data_synch_out => axi_gpio_state
      );
      
    -- AXI control signals from Python
    from_axi.rx_reset      <= axi_gpio_ctrl_async(0); -- async (clk_sys)
    from_axi.tx_reset      <= axi_gpio_ctrl_async(1); -- async (clk_sys)
    from_axi.rx_aligner_en <= axi_gpio_ctrl(2); -- rxusrclk
    from_axi.tx_enc_bypass <= axi_gpio_ctrl(3); -- txusrclk
    -- Rx GT Equalizer
    from_axi.gt_eq.lpmgc   <= axi_gpio_ctrl_async(11 downto 10); -- {gt_ctrl.rxlpmgchold   , gt_ctrl.rxlpmgcovrden  }
    from_axi.gt_eq.lpmhf   <= axi_gpio_ctrl_async( 9 downto  8); -- {gt_ctrl.rxlpmhfhold   , gt_ctrl.rxlpmhfovrden  }
    from_axi.gt_eq.lpmlf   <= axi_gpio_ctrl_async( 7 downto  6); -- {gt_ctrl.rxlpmlfklhold , gt_ctrl.rxlpmlfklovrden}
    from_axi.gt_eq.lpmos   <= axi_gpio_ctrl_async( 5 downto  4); -- {gt_ctrl.rxlpmoshold   , gt_ctrl.rxlpmosovrden  }
    
   bit_synch_axi_to_rx: entity work.bit_synch
    port map (
        bit_in  => axi_gpio_ctrl_async(2), 
        clk     => rxusrclk, 
        bit_out => axi_gpio_ctrl(2)
    ); 
   bit_synch_axi_to_tx: entity work.bit_synch
    port map (
        bit_in  => axi_gpio_ctrl_async(3), 
        clk     => txusrclk, 
        bit_out => axi_gpio_ctrl(3)
    ); 

    ----------------------------------------------------------------------------
    -- UDP to AXI Master
    ----------------------------------------------------------------------------
    
    system_ctrl_inst: entity work.system_control
     port map (

        sys_clk_125 => clk_sys,

        ------------------------------------------------------------------------
        -- 1000 Base-X Transceiver
        ------------------------------------------------------------------------

        -- Ethernet SFP 125 MHz reference clock 
        eth_gtrefclk_p => eth_gtrefclk_p,
        eth_gtrefclk_n => eth_gtrefclk_n,

        -- Ethernet SFP lane
        txn_eth_sfp => txn_eth_sfp,
        txp_eth_sfp => txp_eth_sfp,
        rxn_eth_sfp => rxn_eth_sfp,
        rxp_eth_sfp => rxp_eth_sfp,

        eth_addr_sel   => eth_addr_sel,
        ------------------------------------------------------------------------
        -- I2C Master and GPIOs
        ------------------------------------------------------------------------

        -- I2C Interface (Master)
        sda => sda,
        scl => scl,

        -- DEBUG LEDs
        --GPIO_LED : out std_logic_vector(7 downto 0);

        ------------------------------------------------------------------------
        -- Master AXI-Lite interface
        ------------------------------------------------------------------------

        m_axi_resetn => resetn_axi,

        ---- vectors of AXI Interfaces controlling the Data Lanes
        m_axi_lane_awaddr  => m_axi_lane_awaddr, 
        m_axi_lane_awvalid => m_axi_lane_awvalid,
        m_axi_lane_awready => m_axi_lane_awready,
        m_axi_lane_wdata   => m_axi_lane_wdata,  
        m_axi_lane_wstrb   => m_axi_lane_wstrb,  
        m_axi_lane_wvalid  => m_axi_lane_wvalid, 
        m_axi_lane_wready  => m_axi_lane_wready, 
        m_axi_lane_bresp   => m_axi_lane_bresp,  
        m_axi_lane_bvalid  => m_axi_lane_bvalid, 
        m_axi_lane_bready  => m_axi_lane_bready, 
        m_axi_lane_araddr  => m_axi_lane_araddr, 
        m_axi_lane_arvalid => m_axi_lane_arvalid,
        m_axi_lane_arready => m_axi_lane_arready,
        m_axi_lane_rdata   => m_axi_lane_rdata,  
        m_axi_lane_rresp   => m_axi_lane_rresp,  
        m_axi_lane_rvalid  => m_axi_lane_rvalid, 
        m_axi_lane_rready  => m_axi_lane_rready, 

        ---- Auxiliary Interface
        m_axi_aux_awaddr  => m_axi_aux_awaddr, 
        m_axi_aux_awvalid => m_axi_aux_awvalid,
        m_axi_aux_awready => m_axi_aux_awready,
        m_axi_aux_wdata   => m_axi_aux_wdata,
        m_axi_aux_wstrb   => m_axi_aux_wstrb,  
        m_axi_aux_wvalid  => m_axi_aux_wvalid, 
        m_axi_aux_wready  => m_axi_aux_wready, 
        m_axi_aux_bresp   => m_axi_aux_bresp,  
        m_axi_aux_bvalid  => m_axi_aux_bvalid, 
        m_axi_aux_bready  => m_axi_aux_bready, 
        m_axi_aux_araddr  => m_axi_aux_araddr, 
        m_axi_aux_arvalid => m_axi_aux_arvalid,
        m_axi_aux_arready => m_axi_aux_arready,
        m_axi_aux_rdata   => m_axi_aux_rdata,  
        m_axi_aux_rresp   => m_axi_aux_rresp,  
        m_axi_aux_rvalid  => m_axi_aux_rvalid, 
        m_axi_aux_rready  => m_axi_aux_rready

    );
        
     gpio_axi: entity work.axi_gpio_0  -- Address: 0xFFFF0000
      PORT MAP (
          s_axi_aclk    => clk_sys,
          s_axi_aresetn => resetn_axi,
          s_axi_awaddr  => m_axi_aux_awaddr(8 downto 0),
          s_axi_awvalid => m_axi_aux_awvalid,
          s_axi_awready => m_axi_aux_awready,
          s_axi_wdata   => m_axi_aux_wdata,
          s_axi_wstrb   => m_axi_aux_wstrb,
          s_axi_wvalid  => m_axi_aux_wvalid,
          s_axi_wready  => m_axi_aux_wready,
          s_axi_bresp   => m_axi_aux_bresp,
          s_axi_bvalid  => m_axi_aux_bvalid,
          s_axi_bready  => m_axi_aux_bready,
          s_axi_araddr  => m_axi_aux_araddr(8 downto 0),
          s_axi_arvalid => m_axi_aux_arvalid,
          s_axi_arready => m_axi_aux_arready,
          s_axi_rdata   => m_axi_aux_rdata,
          s_axi_rresp   => m_axi_aux_rresp,
          s_axi_rvalid  => m_axi_aux_rvalid,
          s_axi_rready  => m_axi_aux_rready,
          gpio_io_o     => axi_gpio_ctrl_async,
          gpio2_io_i    => axi_gpio_state
      );
      
     gpio_axi_ddmtd: entity work.axi_gpio_0  -- Address: 0x00000000
      PORT MAP (
          s_axi_aclk    => clk_sys,
          s_axi_aresetn => resetn_axi,
          s_axi_awaddr  => m_axi_lane_awaddr(0)(8 downto 0),
          s_axi_awvalid => m_axi_lane_awvalid(0),
          s_axi_awready => m_axi_lane_awready(0),
          s_axi_wdata   => m_axi_lane_wdata(0),
          s_axi_wstrb   => m_axi_lane_wstrb(0),
          s_axi_wvalid  => m_axi_lane_wvalid(0),
          s_axi_wready  => m_axi_lane_wready(0),
          s_axi_bresp   => m_axi_lane_bresp(0),
          s_axi_bvalid  => m_axi_lane_bvalid(0),
          s_axi_bready  => m_axi_lane_bready(0),
          s_axi_araddr  => m_axi_lane_araddr(0)(8 downto 0),
          s_axi_arvalid => m_axi_lane_arvalid(0),
          s_axi_arready => m_axi_lane_arready(0),
          s_axi_rdata   => m_axi_lane_rdata(0),
          s_axi_rresp   => m_axi_lane_rresp(0),
          s_axi_rvalid  => m_axi_lane_rvalid(0),
          s_axi_rready  => m_axi_lane_rready(0),
          gpio_io_o     => open,
          gpio2_io_i    => to_axi.ddmtd_phase
      );
      
   ila_sys_i: entity work.ila_sys
     PORT MAP (
         clk => clk_sys,
         probe0 => axi_gpio_state,
         probe1 => axi_gpio_ctrl_async
     );
      
--ila_axi : entity work.ila_2
-- PORT MAP (
--	clk => clk_sys,
--	---- WREADY
--	probe0(0) => m_axi_awready, 
--	---- AWADDR
--	probe1 => m_axi_awaddr, 
--	---- BRESP
--	probe2 => m_axi_bresp, 
--	---- BVALID
--	probe3(0) => m_axi_bvalid, 
--	---- BREADY
--	probe4(0) => m_axi_bready, 
--	---- ARADDR
--	probe5 => m_axi_araddr, 
--	---- RREADY
--	probe6(0) => m_axi_rready, 
--	---- WVALID
--	probe7(0) => m_axi_wvalid, 
--	---- ARVALID
--	probe8(0) => m_axi_arvalid, 
--	---- ARREADY
--	probe9(0) => m_axi_arready, 
--	---- RDATA
--	probe10 => m_axi_rdata, 
--	---- AWVALID
--	probe11(0) => m_axi_awvalid, 
--	---- AWREADY
--	probe12(0) => m_axi_awready, 
--	---- RRESP
--	probe13 => m_axi_rresp, 
--	---- WDATA
--	probe14 => m_axi_wdata, 
--	---- WSTRB
--	probe15 => m_axi_wstrb, 
--	---- RVALID
--	probe16(0) => m_axi_rvalid, 
--	---- ARPROT
--	probe17 => (others => '0'),
--	---- AWPROT 
--	probe18 => (others => '0') 
--);


end Behavioral;
